module phase_detector
(
input clk,
input a,
input b,
output logic c
);



endmodule
