module half_matrix_dot_vector
#(
parameter WIDTH = 10,
parameter HEIGHT = 10
)
(
input clk,

);

endmodule
